VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_vsdnand4_1x
  CLASS CORE ;
  FOREIGN sky130_vsdnand4_1x ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.970 0.990 2.210 1.660 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.140 0.990 1.450 1.320 ;
        RECT 1.140 0.820 1.350 0.990 ;
        RECT 1.000 0.300 1.350 0.820 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.590 0.990 0.970 1.320 ;
        RECT 0.590 0.300 0.810 0.990 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.990 0.390 1.320 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.080 0.080 0.420 0.820 ;
        RECT 0.000 -0.090 2.300 0.080 ;
      LAYER mcon ;
        RECT 0.140 -0.090 0.310 0.080 ;
        RECT 0.600 -0.090 0.770 0.080 ;
        RECT 1.060 -0.090 1.230 0.080 ;
        RECT 1.520 -0.090 1.690 0.080 ;
        RECT 1.980 -0.090 2.150 0.080 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 -0.090 0.320 0.080 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.300 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.300 2.800 ;
        RECT 0.080 2.480 0.340 2.630 ;
        RECT 0.080 1.490 0.310 2.480 ;
        RECT 1.010 1.830 1.210 2.630 ;
        RECT 1.910 1.830 2.190 2.630 ;
      LAYER mcon ;
        RECT 0.140 2.630 0.310 2.800 ;
        RECT 0.600 2.630 0.770 2.800 ;
        RECT 1.060 2.630 1.230 2.800 ;
        RECT 1.520 2.630 1.690 2.800 ;
        RECT 1.980 2.630 2.150 2.800 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 0.510 1.660 0.840 2.460 ;
        RECT 1.380 1.660 1.710 2.460 ;
        RECT 0.510 1.490 1.790 1.660 ;
        RECT 1.620 0.820 1.790 1.490 ;
        RECT 1.520 0.250 2.210 0.820 ;
    END
  END Y
END sky130_vsdnand4_1x
END LIBRARY

