magic
tech sky130A
timestamp 1615482986
<< nwell >>
rect -19 130 203 291
<< pwell >>
rect 15 -9 32 8
<< nmos >>
rect 39 23 55 88
rect 81 23 96 88
rect 129 23 144 88
<< pmos >>
rect 39 148 55 248
rect 84 148 99 248
rect 129 148 144 248
<< ndiff >>
rect 11 49 39 88
rect 11 32 15 49
rect 32 32 39 49
rect 11 23 39 32
rect 55 23 81 88
rect 96 23 129 88
rect 144 85 171 88
rect 144 84 175 85
rect 144 67 150 84
rect 167 67 175 84
rect 144 50 175 67
rect 144 33 150 50
rect 167 33 175 50
rect 144 25 175 33
rect 144 23 171 25
<< pdiff >>
rect 1 242 39 248
rect 1 225 13 242
rect 30 225 39 242
rect 1 208 39 225
rect 1 191 13 208
rect 30 191 39 208
rect 1 174 39 191
rect 1 157 12 174
rect 29 157 39 174
rect 1 148 39 157
rect 55 238 84 248
rect 55 221 61 238
rect 78 221 84 238
rect 55 204 84 221
rect 55 187 61 204
rect 78 187 84 204
rect 55 170 84 187
rect 55 153 61 170
rect 78 153 84 170
rect 55 148 84 153
rect 99 242 129 248
rect 99 225 105 242
rect 122 225 129 242
rect 99 208 129 225
rect 99 191 105 208
rect 122 191 129 208
rect 99 148 129 191
rect 144 246 173 248
rect 144 242 175 246
rect 144 225 150 242
rect 167 225 175 242
rect 144 208 175 225
rect 144 191 150 208
rect 167 191 175 208
rect 144 174 175 191
rect 144 157 150 174
rect 167 157 175 174
rect 144 149 175 157
rect 144 148 173 149
<< ndiffc >>
rect 15 32 32 49
rect 150 67 167 84
rect 150 33 167 50
<< pdiffc >>
rect 13 225 30 242
rect 13 191 30 208
rect 12 157 29 174
rect 61 221 78 238
rect 61 187 78 204
rect 61 153 78 170
rect 105 225 122 242
rect 105 191 122 208
rect 150 225 167 242
rect 150 191 167 208
rect 150 157 167 174
<< poly >>
rect 39 248 55 261
rect 84 248 99 261
rect 129 248 144 261
rect 39 132 55 148
rect 11 124 55 132
rect 84 132 99 148
rect 129 132 144 148
rect 84 130 108 132
rect 11 107 16 124
rect 33 107 55 124
rect 11 99 55 107
rect 39 88 55 99
rect 81 124 108 130
rect 81 107 86 124
rect 103 107 108 124
rect 81 99 108 107
rect 129 124 175 132
rect 129 107 147 124
rect 164 107 175 124
rect 129 102 175 107
rect 81 88 96 99
rect 129 88 144 102
rect 39 10 55 23
rect 81 10 96 23
rect 129 10 144 23
<< polycont >>
rect 16 107 33 124
rect 86 107 103 124
rect 147 107 164 124
<< locali >>
rect 0 263 14 280
rect 31 263 60 280
rect 77 263 106 280
rect 123 263 152 280
rect 169 263 184 280
rect 9 242 34 263
rect 9 225 13 242
rect 30 225 34 242
rect 9 208 34 225
rect 9 191 13 208
rect 30 191 34 208
rect 9 174 34 191
rect 9 157 12 174
rect 29 157 34 174
rect 9 149 34 157
rect 51 238 84 246
rect 51 221 61 238
rect 78 221 84 238
rect 51 204 84 221
rect 51 187 61 204
rect 78 187 84 204
rect 51 170 84 187
rect 101 242 124 263
rect 101 225 105 242
rect 122 225 124 242
rect 101 208 124 225
rect 101 191 105 208
rect 122 191 124 208
rect 101 183 124 191
rect 141 242 175 246
rect 141 225 150 242
rect 167 225 175 242
rect 141 208 175 225
rect 141 191 150 208
rect 167 191 175 208
rect 51 153 61 170
rect 78 166 84 170
rect 141 174 175 191
rect 141 166 150 174
rect 78 157 150 166
rect 167 157 175 174
rect 78 153 175 157
rect 51 149 175 153
rect 11 124 33 132
rect 11 107 16 124
rect 11 74 33 107
rect 51 59 69 149
rect 86 124 122 132
rect 103 107 122 124
rect 86 76 122 107
rect 139 124 175 132
rect 139 107 147 124
rect 164 107 175 124
rect 139 102 175 107
rect 141 84 175 85
rect 141 67 150 84
rect 167 67 175 84
rect 141 59 175 67
rect 9 49 34 57
rect 9 32 15 49
rect 32 32 34 49
rect 9 8 34 32
rect 51 50 175 59
rect 51 33 150 50
rect 167 33 175 50
rect 51 25 175 33
rect 0 -9 14 8
rect 31 -9 60 8
rect 77 -9 106 8
rect 123 -9 152 8
rect 169 -9 184 8
<< viali >>
rect 14 263 31 280
rect 60 263 77 280
rect 106 263 123 280
rect 152 263 169 280
rect 14 -9 31 8
rect 60 -9 77 8
rect 106 -9 123 8
rect 152 -9 169 8
<< metal1 >>
rect 0 280 184 296
rect 0 263 14 280
rect 31 263 60 280
rect 77 263 106 280
rect 123 263 152 280
rect 169 263 184 280
rect 0 248 184 263
rect 0 8 184 24
rect 0 -9 14 8
rect 31 -9 60 8
rect 77 -9 106 8
rect 123 -9 152 8
rect 169 -9 184 8
rect 0 -24 184 -9
<< labels >>
flabel locali s 61 42 78 59 0 FreeSans 125 0 0 0 Y
port 8 nsew signal output
flabel locali s 153 110 170 127 0 FreeSans 125 0 0 0 A
port 1 nsew signal input
flabel locali s 15 110 32 127 0 FreeSans 125 0 0 0 C
port 3 nsew signal input
flabel locali s 107 110 124 127 0 FreeSans 125 0 0 0 B
port 2 nsew signal input
flabel pwell s 15 -9 32 8 0 FreeSans 100 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 15 -9 32 8 0 FreeSans 100 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 15 263 32 280 0 FreeSans 100 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand3_1
flabel nwell s 15 263 32 280 0 FreeSans 100 0 0 0 VPB
port 6 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite unithd
string FIXED_BBOX 0 0 184 272
string LEFsymmetry X Y R90
string path 0.000 0.000 9.200 0.000 
<< end >>
