VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_vsdnand3_1x
  CLASS CORE ;
  FOREIGN sky130_vsdnand3_1x ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.390 1.020 1.750 1.320 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.860 0.760 1.220 1.320 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.264000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.740 0.330 1.320 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.080 0.340 0.570 ;
        RECT 0.000 -0.090 1.840 0.080 ;
      LAYER mcon ;
        RECT 0.140 -0.090 0.310 0.080 ;
        RECT 0.600 -0.090 0.770 0.080 ;
        RECT 1.060 -0.090 1.230 0.080 ;
        RECT 1.520 -0.090 1.690 0.080 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 -0.090 0.320 0.080 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.300 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.800 ;
        RECT 0.090 1.490 0.340 2.630 ;
        RECT 1.010 1.830 1.240 2.630 ;
      LAYER mcon ;
        RECT 0.140 2.630 0.310 2.800 ;
        RECT 0.600 2.630 0.770 2.800 ;
        RECT 1.060 2.630 1.230 2.800 ;
        RECT 1.520 2.630 1.690 2.800 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.798900 ;
    PORT
      LAYER li1 ;
        RECT 0.510 1.660 0.840 2.460 ;
        RECT 1.410 1.660 1.750 2.460 ;
        RECT 0.510 1.490 1.750 1.660 ;
        RECT 0.510 0.590 0.690 1.490 ;
        RECT 1.410 0.590 1.750 0.850 ;
        RECT 0.510 0.250 1.750 0.590 ;
    END
  END Y
END sky130_vsdnand3_1x
END LIBRARY

