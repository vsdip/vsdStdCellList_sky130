* SPICE3 file created from sky130_vsdinv_8x.ext - technology: sky130A

.option scale=0.01u

.subckt sky130_vsdinv_8x A Y VPWR VGND VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=66 l=15
X1 VGND A Y VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=66 l=15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=66 l=15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=66 l=15
X5 Y A VGND VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X6 VGND A Y VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X7 Y A VGND VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X8 VGND A Y VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X9 VGND A Y VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=66 l=15
X11 Y A VGND VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=66 l=15
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=66 l=15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=66 l=15
X15 Y A VGND VGND sky130_fd_pr__nfet_01v8 w=42 l=15

.ends
