* SPICE3 file created from sky130_vsd_conb.ext - technology: sky130A

.option scale=10000u

.subckt sky130_vsd_conb HI LO VGND VPB
X0 VPB LO HI w_n13_156# sky130_fd_pr__pfet_01v8 w=60 l=15
X1 HI HI VPB w_n13_156# sky130_fd_pr__pfet_01v8 w=60 l=15
X2 LO HI VGND VGND sky130_fd_pr__nfet_01v8 w=42 l=15
X3 VGND LO LO VGND sky130_fd_pr__nfet_01v8 w=42 l=15
C0 HI LO 0.13fF
C1 w_n13_156# VPB 0.02fF
C2 w_n13_156# HI 0.00fF
C3 LO VPB 0.03fF
C4 HI VPB 0.16fF
C5 VPB VGND 0.30fF
C6 LO VGND 0.33fF
C7 HI VGND 0.32fF
C8 w_n13_156# VGND 0.27fF
.ends
