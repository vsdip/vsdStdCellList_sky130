VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_vsdclkbuf_4x
  CLASS CORE ;
  FOREIGN sky130_vsdclkbuf_4x ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.214500 ;
    PORT
      LAYER li1 ;
        RECT 0.420 0.780 0.770 1.320 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.943800 ;
    PORT
      LAYER li1 ;
        RECT 1.050 2.000 1.310 2.460 ;
        RECT 1.980 2.000 2.320 2.460 ;
        RECT 1.050 1.830 2.320 2.000 ;
        RECT 1.980 1.580 2.320 1.830 ;
        RECT 1.980 1.410 2.820 1.580 ;
        RECT 2.410 0.980 2.820 1.410 ;
        RECT 2.320 0.910 2.820 0.980 ;
        RECT 2.150 0.900 2.820 0.910 ;
        RECT 1.020 0.800 2.820 0.900 ;
        RECT 1.020 0.740 2.490 0.800 ;
        RECT 1.020 0.730 2.320 0.740 ;
        RECT 1.020 0.340 1.310 0.730 ;
        RECT 1.990 0.280 2.320 0.730 ;
    END
  END Y
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.920 2.800 ;
        RECT 0.560 1.830 0.880 2.630 ;
        RECT 1.500 2.170 1.760 2.630 ;
        RECT 2.490 1.760 2.780 2.630 ;
      LAYER mcon ;
        RECT 0.140 2.630 0.310 2.800 ;
        RECT 0.600 2.630 0.770 2.800 ;
        RECT 1.070 2.630 1.240 2.800 ;
        RECT 1.550 2.630 1.720 2.800 ;
        RECT 2.060 2.630 2.230 2.800 ;
        RECT 2.600 2.630 2.770 2.800 ;
      LAYER met1 ;
        RECT 0.000 2.550 2.920 2.960 ;
    END
  END VPWR
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.300 3.110 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140 -0.090 0.310 0.080 ;
      LAYER li1 ;
        RECT 0.550 0.080 0.830 0.570 ;
        RECT 1.490 0.280 1.820 0.560 ;
        RECT 1.500 0.080 1.760 0.280 ;
        RECT 2.490 0.080 2.770 0.570 ;
        RECT 0.000 -0.170 2.920 0.080 ;
      LAYER mcon ;
        RECT 0.140 -0.090 0.310 0.080 ;
        RECT 0.600 -0.090 0.770 0.080 ;
        RECT 1.070 -0.090 1.240 0.080 ;
        RECT 1.550 -0.090 1.720 0.080 ;
        RECT 2.060 -0.090 2.230 0.080 ;
        RECT 2.600 -0.090 2.770 0.080 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.920 0.180 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.080 1.660 0.390 2.460 ;
        RECT 0.080 1.490 1.120 1.660 ;
        RECT 0.080 0.590 0.250 1.490 ;
        RECT 0.940 1.240 1.120 1.490 ;
        RECT 0.940 1.070 1.980 1.240 ;
        RECT 0.080 0.250 0.380 0.590 ;
  END
END sky130_vsdclkbuf_4x
END LIBRARY

