VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_vsdo21ai_1x
  CLASS CORE ;
  FOREIGN sky130_vsdo21ai_1x ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.080 0.950 0.410 1.610 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.600 1.340 0.770 1.640 ;
        RECT 0.600 1.040 1.000 1.340 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.510 1.350 1.730 1.680 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.550 0.080 0.880 0.440 ;
        RECT 0.000 -0.090 1.840 0.080 ;
      LAYER mcon ;
        RECT 0.140 -0.090 0.310 0.080 ;
        RECT 0.600 -0.090 0.770 0.080 ;
        RECT 1.060 -0.090 1.230 0.080 ;
        RECT 1.520 -0.090 1.690 0.080 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140 -0.090 0.310 0.080 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.300 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.800 ;
        RECT 0.140 1.820 0.470 2.630 ;
        RECT 1.470 1.850 1.720 2.630 ;
      LAYER mcon ;
        RECT 0.140 2.630 0.310 2.800 ;
        RECT 0.600 2.630 0.770 2.800 ;
        RECT 1.060 2.630 1.230 2.800 ;
        RECT 1.520 2.630 1.690 2.800 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299000 ;
    PORT
      LAYER li1 ;
        RECT 0.960 1.680 1.300 2.460 ;
        RECT 0.960 1.510 1.340 1.680 ;
        RECT 1.170 1.120 1.340 1.510 ;
        RECT 1.170 0.950 1.740 1.120 ;
        RECT 1.450 0.280 1.740 0.950 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.120 0.610 1.280 0.780 ;
        RECT 0.120 0.280 0.380 0.610 ;
        RECT 1.050 0.280 1.280 0.610 ;
  END
END sky130_vsdo21ai_1x
END LIBRARY

