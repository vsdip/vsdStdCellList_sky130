magic
tech sky130A
timestamp 1616139194
<< nwell >>
rect -8 160 436 292
rect 18 159 424 160
<< nmos >>
rect 46 38 61 80
rect 90 38 105 80
rect 137 38 152 80
rect 183 38 198 80
rect 230 38 245 80
rect 277 38 292 80
rect 326 38 341 80
rect 373 38 388 80
<< pmos >>
rect 46 180 61 246
rect 90 180 105 246
rect 137 180 152 246
rect 183 180 198 246
rect 230 180 245 246
rect 277 180 292 246
rect 326 180 341 246
rect 373 180 388 246
<< ndiff >>
rect 18 63 46 80
rect 18 46 22 63
rect 39 46 46 63
rect 18 38 46 46
rect 61 64 90 80
rect 61 47 67 64
rect 84 47 90 64
rect 61 38 90 47
rect 105 60 137 80
rect 105 43 114 60
rect 131 43 137 60
rect 105 38 137 43
rect 152 65 183 80
rect 152 48 159 65
rect 176 48 183 65
rect 152 38 183 48
rect 198 60 230 80
rect 198 43 206 60
rect 223 43 230 60
rect 198 38 230 43
rect 245 65 277 80
rect 245 48 254 65
rect 271 48 277 65
rect 245 38 277 48
rect 292 60 326 80
rect 292 43 300 60
rect 317 43 326 60
rect 292 38 326 43
rect 341 65 373 80
rect 341 48 349 65
rect 366 48 373 65
rect 341 38 373 48
rect 388 59 422 80
rect 388 42 398 59
rect 415 42 422 59
rect 388 38 422 42
<< pdiff >>
rect 20 246 37 257
rect 15 239 46 246
rect 15 206 20 239
rect 37 206 46 239
rect 15 180 46 206
rect 61 232 90 246
rect 61 194 67 232
rect 84 194 90 232
rect 61 180 90 194
rect 105 240 137 246
rect 105 203 112 240
rect 129 203 137 240
rect 105 180 137 203
rect 152 232 183 246
rect 152 186 159 232
rect 176 186 183 232
rect 152 180 183 186
rect 198 239 230 246
rect 198 199 205 239
rect 222 199 230 239
rect 198 180 230 199
rect 245 231 277 246
rect 245 190 253 231
rect 270 190 277 231
rect 245 180 277 190
rect 292 240 326 246
rect 292 199 300 240
rect 317 199 326 240
rect 292 180 326 199
rect 341 233 373 246
rect 341 192 349 233
rect 366 192 373 233
rect 341 180 373 192
rect 388 240 418 246
rect 388 199 397 240
rect 414 199 418 240
rect 388 180 418 199
<< ndiffc >>
rect 22 46 39 63
rect 67 47 84 64
rect 114 43 131 60
rect 159 48 176 65
rect 206 43 223 60
rect 254 48 271 65
rect 300 43 317 60
rect 349 48 366 65
rect 398 42 415 59
<< pdiffc >>
rect 20 206 37 239
rect 67 194 84 232
rect 112 203 129 240
rect 159 186 176 232
rect 205 199 222 239
rect 253 190 270 231
rect 300 199 317 240
rect 349 192 366 233
rect 397 199 414 240
<< psubdiff >>
rect 3 9 420 11
rect 3 -8 45 9
rect 62 -8 87 9
rect 104 -8 129 9
rect 146 -8 172 9
rect 189 -8 216 9
rect 233 -8 258 9
rect 275 -8 301 9
rect 318 -8 347 9
rect 364 -8 420 9
<< psubdiffcont >>
rect 45 -8 62 9
rect 87 -8 104 9
rect 129 -8 146 9
rect 172 -8 189 9
rect 216 -8 233 9
rect 258 -8 275 9
rect 301 -8 318 9
rect 347 -8 364 9
<< poly >>
rect 46 246 61 259
rect 90 246 105 259
rect 137 246 152 259
rect 183 246 198 259
rect 230 246 245 259
rect 277 246 292 259
rect 326 246 341 260
rect 373 246 388 260
rect 46 141 61 180
rect 90 141 105 180
rect 137 141 152 180
rect 183 141 198 180
rect 230 141 245 180
rect 277 141 292 180
rect 326 141 341 180
rect 373 141 388 180
rect 38 136 388 141
rect 38 119 46 136
rect 63 119 80 136
rect 97 119 114 136
rect 131 119 148 136
rect 165 119 182 136
rect 199 119 217 136
rect 234 119 251 136
rect 268 119 285 136
rect 302 119 319 136
rect 336 119 353 136
rect 370 119 388 136
rect 38 114 388 119
rect 46 80 61 114
rect 90 80 105 114
rect 137 80 152 114
rect 183 80 198 114
rect 230 80 245 114
rect 277 80 292 114
rect 326 80 341 114
rect 373 80 388 114
rect 46 23 61 38
rect 90 23 105 38
rect 137 23 152 38
rect 183 23 198 38
rect 230 23 245 38
rect 277 23 292 38
rect 326 24 341 38
rect 373 24 388 38
<< polycont >>
rect 46 119 63 136
rect 80 119 97 136
rect 114 119 131 136
rect 148 119 165 136
rect 182 119 199 136
rect 217 119 234 136
rect 251 119 268 136
rect 285 119 302 136
rect 319 119 336 136
rect 353 119 370 136
<< locali >>
rect 2 280 422 282
rect 2 263 4 280
rect 21 263 46 280
rect 63 263 84 280
rect 101 263 129 280
rect 146 263 171 280
rect 188 263 216 280
rect 233 263 255 280
rect 272 279 397 280
rect 272 263 301 279
rect 2 262 301 263
rect 318 262 348 279
rect 365 263 397 279
rect 414 263 422 280
rect 365 262 422 263
rect 2 261 422 262
rect 20 239 37 261
rect 20 191 37 206
rect 67 232 84 241
rect 67 174 84 194
rect 112 240 129 261
rect 112 191 129 203
rect 159 232 176 241
rect 205 239 222 261
rect 205 191 222 199
rect 253 231 270 241
rect 159 174 176 186
rect 300 240 317 261
rect 300 191 317 199
rect 349 233 366 241
rect 253 174 270 190
rect 349 174 366 192
rect 397 240 414 261
rect 397 191 414 199
rect 0 154 426 174
rect 0 98 21 154
rect 38 136 391 137
rect 38 119 46 136
rect 63 119 80 136
rect 97 119 114 136
rect 131 119 148 136
rect 165 119 182 136
rect 199 119 217 136
rect 234 119 251 136
rect 268 119 285 136
rect 302 119 319 136
rect 336 119 353 136
rect 370 119 391 136
rect 409 98 426 154
rect 0 81 426 98
rect 66 80 426 81
rect 67 64 84 80
rect 14 63 48 64
rect 14 46 22 63
rect 39 46 48 63
rect 14 39 48 46
rect 159 65 176 80
rect 14 38 43 39
rect 67 38 84 47
rect 104 60 139 63
rect 104 43 114 60
rect 131 43 139 60
rect 104 38 139 43
rect 254 65 271 80
rect 159 38 176 48
rect 198 60 231 63
rect 198 43 206 60
rect 223 43 231 60
rect 198 38 231 43
rect 349 65 366 80
rect 254 38 271 48
rect 292 60 325 63
rect 292 43 300 60
rect 317 43 325 60
rect 20 11 37 38
rect 3 10 37 11
rect 114 10 131 38
rect 206 10 223 38
rect 300 10 317 43
rect 349 38 366 48
rect 390 59 423 62
rect 390 42 398 59
rect 415 42 423 59
rect 390 38 423 42
rect 396 10 413 38
rect 3 9 421 10
rect 20 -8 45 9
rect 62 -8 87 9
rect 104 -8 129 9
rect 146 -8 172 9
rect 189 -8 216 9
rect 233 -8 258 9
rect 275 -8 301 9
rect 318 -8 347 9
rect 364 -8 396 9
rect 413 -8 421 9
rect 3 -10 421 -8
<< viali >>
rect 4 263 21 280
rect 46 263 63 280
rect 84 263 101 280
rect 129 263 146 280
rect 171 263 188 280
rect 216 263 233 280
rect 255 263 272 280
rect 301 262 318 279
rect 348 262 365 279
rect 397 263 414 280
rect 3 -8 20 9
rect 45 -8 62 9
rect 87 -8 104 9
rect 129 -8 146 9
rect 172 -8 189 9
rect 216 -8 233 9
rect 258 -8 275 9
rect 301 -8 318 9
rect 347 -8 364 9
rect 396 -8 413 9
<< metal1 >>
rect 0 280 428 290
rect 0 263 4 280
rect 21 263 46 280
rect 63 263 84 280
rect 101 263 129 280
rect 146 263 171 280
rect 188 263 216 280
rect 233 263 255 280
rect 272 279 397 280
rect 272 263 301 279
rect 0 262 301 263
rect 318 262 348 279
rect 365 263 397 279
rect 414 263 428 280
rect 365 262 428 263
rect 0 252 428 262
rect 20 191 37 252
rect 0 9 428 19
rect 0 -8 3 9
rect 20 -8 45 9
rect 62 -8 87 9
rect 104 -8 129 9
rect 146 -8 172 9
rect 189 -8 216 9
rect 233 -8 258 9
rect 275 -8 301 9
rect 318 -8 347 9
rect 364 -8 396 9
rect 413 -8 428 9
rect 0 -20 428 -8
<< labels >>
flabel metal1 189 -10 216 10 0 FreeSans 120 0 0 0 VGND
port 4 nsew ground bidirectional
flabel nwell 4 263 21 280 0 FreeSans 1 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 188 261 216 282 0 FreeSans 120 0 0 0 VPWR
port 3 nsew power bidirectional
flabel locali 370 119 391 137 0 FreeSans 120 0 0 0 A
port 1 nsew signal input
flabel locali 409 80 426 174 0 FreeSans 120 0 0 0 Y
port 2 nsew signal output
<< properties >>
string LEFclass CORE
string LEFsite unithd
string FIXED_BBOX 0 0 428 272
string LEFsymmetry X Y R90
<< end >>
